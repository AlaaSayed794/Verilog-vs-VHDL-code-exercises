module Switches_to_LEDs (
    input i1,
    input i2,
    input i3,
    output o1,
    output o2,
    output o3
);
assign o1 = i1;
assign o2 = i2;
assign o3 = i3;    
endmodule