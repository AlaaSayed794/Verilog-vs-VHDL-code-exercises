module AND_gate (
    input i1,
    input i2,
    output o1
);
assign o1 = i1 & i2; 
endmodule