library ieee;
use ieee.std_logic_1164.all ;

entity AND_gate is 
port(
    i1 : in std_logic;
    i2 : in std_logic;
    o1 : out std_logic;
    );
end entity AND_gate;

architecture RTL of AND_gate is
    begin
        o1 <= i1 and i2;
end architecture RTL;